// +FHDR============================================================================/
// Author       : huangjie
// Creat Time   : 2023/06/19 14:12:50
// File Name    : iic_m_phy_warper.v
// Module Ver   : Vx.x
//
//
// All Rights Reserved
//
// ---------------------------------------------------------------------------------/
//
// Modification History:
// V1.0         initial
//
// -FHDR============================================================================/
// 
// iic_m_phy_warper
//    |---
// 
`timescale 1ns/1ps

module iic_m_phy_warper #
(
    parameter                           U_DLY = 1                     // 
)
(
// ---------------------------------------------------------------------------------
// CLock & Reset
// ---------------------------------------------------------------------------------
    input                               clk_sys                     ,
    input                               rst_n                       ,
// ---------------------------------------------------------------------------------
// Config
// ---------------------------------------------------------------------------------
    input                               baud_en                     , 
// ---------------------------------------------------------------------------------
// User Data
// ---------------------------------------------------------------------------------
    output                              usr_wready                  , 
    input                               usr_wvalid                  , 
    input                         [3:0] usr_wcmd                    , // bit3 -> master ack status,bit2 -> rd/wrn,bit1 -> end,bit0->start.
    input                         [7:0] usr_wdata                   , 

    output                        [7:0] usr_rdata                   , 
    output                              usr_rvalid                  , 
// ---------------------------------------------------------------------------------
// IIC Phy
// ---------------------------------------------------------------------------------
    input                               iic_sck_i                   , 
    output                              iic_sck_o                   , 
    output                              iic_sck_t                   , 
    input                               iic_sda_i                   , 
    output                              iic_sda_o                   , 
    output                              iic_sda_t                   , 
// ---------------------------------------------------------------------------------
// Debug
// ---------------------------------------------------------------------------------
    output                              dgb_err_sack                , 
    output                              dbg_err_abt                   
);

wire                                    bit_wready                  ; 
wire                                    bit_wvalid                  ; 
wire                             [11:0] bit_wdata                   ; 

wire                                    bit_rdata                   ; 
wire                                    bit_rvalid                  ; 

iic_m_phy_bitgen #
(
    .U_DLY                          (U_DLY                      )  // 
)
u_iic_m_phy_bitgen
(
// ---------------------------------------------------------------------------------
// CLock & Reset
// ---------------------------------------------------------------------------------
    .clk_sys                        (clk_sys                    ), // (input )
    .rst_n                          (rst_n                      ), // (input )
// ---------------------------------------------------------------------------------
// User Data
// ---------------------------------------------------------------------------------
    .usr_wready                     (usr_wready                 ), // (output)
    .usr_wvalid                     (usr_wvalid                 ), // (input )
    .usr_wcmd                       (usr_wcmd[3:0]              ), // (input ) bit3 -> master ack status,bit2 -> rd/wrn,bit1 -> end,bit0->start.
    .usr_wdata                      (usr_wdata[7:0]             ), // (input )

    .usr_rdata                      (usr_rdata[7:0]             ), // (output)
    .usr_rvalid                     (usr_rvalid                 ), // (output)
// ---------------------------------------------------------------------------------
// Bit Data
// ---------------------------------------------------------------------------------
    .bit_wready                     (bit_wready                 ), // (input )
    .bit_wvalid                     (bit_wvalid                 ), // (output)
    .bit_wdata                      (bit_wdata[11:0]            ), // (output)

    .bit_rdata                      (bit_rdata                  ), // (input )
    .bit_rvalid                     (bit_rvalid                 ), // (input )
// ---------------------------------------------------------------------------------
// Debug
// ---------------------------------------------------------------------------------
    .dgb_err_sack                   (dgb_err_sack               )  // (output)
);

iic_m_phy_timing #
(
    .U_DLY                          (U_DLY                      )  // 
)
u_iic_m_phy_timing
(
// ---------------------------------------------------------------------------------
// CLock & Reset
// ---------------------------------------------------------------------------------
    .clk_sys                        (clk_sys                    ), // (input )
    .rst_n                          (rst_n                      ), // (input )
// ---------------------------------------------------------------------------------
// Baud
// ---------------------------------------------------------------------------------
    .baud_en                        (baud_en                    ), // (input )
// ---------------------------------------------------------------------------------
// Bit Data
// ---------------------------------------------------------------------------------
    .bit_wready                     (bit_wready                 ), // (output)
    .bit_wvalid                     (bit_wvalid                 ), // (input )
    .bit_wdata                      (bit_wdata[11:0]            ), // (input )

    .bit_rdata                      (bit_rdata                  ), // (output)
    .bit_rvalid                     (bit_rvalid                 ), // (output)
// ---------------------------------------------------------------------------------
// IIC Phy
// ---------------------------------------------------------------------------------
    .iic_sck_i                      (iic_sck_i                  ), // (input )
    .iic_sck_o                      (iic_sck_o                  ), // (output)
    .iic_sck_t                      (iic_sck_t                  ), // (output)
    .iic_sda_i                      (iic_sda_i                  ), // (input )
    .iic_sda_o                      (iic_sda_o                  ), // (output)
    .iic_sda_t                      (iic_sda_t                  ), // (output)
// ---------------------------------------------------------------------------------
// Debug
// ---------------------------------------------------------------------------------
    .dbg_err_abt                    (dbg_err_abt                )  // (output)
);

endmodule

